package types;
    typedef enum bit [1:0] {DS1, PS, SS, DS0} sreg_index_e;
endpackage
